library ieee;
use ieee.std_logic_1164.all;

entity FF_tipoT is
	port(clk: in std_logic;
			q : buffer std_logic);
end FF_tipoT;

architecture arc_FF_TipoT of FF_tipoT is
	signal s: std_logic;
begin
	s <= q;
	process(clk)
	begin
		if clk'event and clk = '1' then
			s <= not s;
		end if;
		q <= s;
	end process;
end arc_FF_TipoT;